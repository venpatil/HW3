/////////////////////////////////////////////
// Simple SystemVerilog Package
// ece571_cpu_pkg.sv
// Makes use of parameter, enum, and struct
// Venkatesh Patil (venpatil@pdx.edu)
// Modify to add your content
////////////////////////////////////////////

package ece571_cpu_pkg;

// Parameter for ALU size



// Enumeration for opcodes




// Packed structs for instructions



endpackage
