////////////////////////////////////////////////
// Simple 5-stage pipelined CPU
//  But we will not use the Memory/Regfile
// It will only be for connectivity
// // ece571_cpu.sv
// Venkatesh Patil (venpatil@pdx.edu)
// Modify as needed
// For ECE571 hw3 labs use
///////////////////////////////////////////////

module ece571_cpu (

  //ports declarations 

   //Piplined Registers


  // Instantiate modules

  // Pipelining Logic
 


endmodule
