//////////////////////////////////////////////
// Simple ALU operations 
// Venkatesh patil (venpatil@pdx.edu
// To be used with ECE-571 HW3 labs
// Modify as needed
// 
// Make use of package to get the opcodes

////////////////////////////////////////////

// ece571_alu.sv
module ece571_alu (



endmodule
